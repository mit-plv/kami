import Vector::*;
import BuildVector::*;
import RegFile::*;
import RegFileZero::*;
import FIFO::*;
import FIFOF::*;
import SimpleBRAM::*;
import MulDiv::*;
import SpecialFIFOs::*;


