// The CC interface is defined in the header part (thus in Header.bsv)
