interface Mem;
    method Action mem_enq_rq_0 (Struct2 rq);
    method ActionValue#(Struct2) mem_deq_rs_0 ();
    method Action mem_enq_rq_1 (Struct2 rq);
    method ActionValue#(Struct2) mem_deq_rs_1 ();
    method Action mem_enq_rq_2 (Struct2 rq);
    method ActionValue#(Struct2) mem_deq_rs_2 ();
    method Action mem_enq_rq_3 (Struct2 rq);
    method ActionValue#(Struct2) mem_deq_rs_3 ();
    method Action mem_enq_rq_4 (Struct2 rq);
    method ActionValue#(Struct2) mem_deq_rs_4 ();
    method Action mem_enq_rq_5 (Struct2 rq);
    method ActionValue#(Struct2) mem_deq_rs_5 ();
    method Action mem_enq_rq_6 (Struct2 rq);
    method ActionValue#(Struct2) mem_deq_rs_6 ();
    method Action mem_enq_rq_7 (Struct2 rq);
    method ActionValue#(Struct2) mem_deq_rs_7 ();

    method Bool isInit ();
endinterface
