import Vector::*;
import BuildVector::*;
import RegFile::*;
import FIFO::*;
import FIFOF::*;
import SimpleBRAM::*;
import MulDiv::*;
import SpecialFIFOs::*;

interface Proc;
endinterface

